module BramMem(
  input         clock,
  input  [4:0]  io_addr, // @[\\src\\main\\scala\\bram\\bramMem.scala 32:14]
  input         io_en, // @[\\src\\main\\scala\\bram\\bramMem.scala 32:14]
  input         io_wrEn, // @[\\src\\main\\scala\\bram\\bramMem.scala 32:14]
  input  [27:0] io_wrData, // @[\\src\\main\\scala\\bram\\bramMem.scala 32:14]
  output [27:0] io_rdData // @[\\src\\main\\scala\\bram\\bramMem.scala 32:14]
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [27:0] mem [0:27]; // @[\\src\\main\\scala\\bram\\bramMem.scala 43:24]
  wire  mem_io_rdData_MPORT_en; // @[\\src\\main\\scala\\bram\\bramMem.scala 43:24]
  wire [4:0] mem_io_rdData_MPORT_addr; // @[\\src\\main\\scala\\bram\\bramMem.scala 43:24]
  wire [27:0] mem_io_rdData_MPORT_data; // @[\\src\\main\\scala\\bram\\bramMem.scala 43:24]
  wire [27:0] mem_MPORT_data; // @[\\src\\main\\scala\\bram\\bramMem.scala 43:24]
  wire [4:0] mem_MPORT_addr; // @[\\src\\main\\scala\\bram\\bramMem.scala 43:24]
  wire  mem_MPORT_mask; // @[\\src\\main\\scala\\bram\\bramMem.scala 43:24]
  wire  mem_MPORT_en; // @[\\src\\main\\scala\\bram\\bramMem.scala 43:24]
  reg  mem_io_rdData_MPORT_en_pipe_0;
  reg [4:0] mem_io_rdData_MPORT_addr_pipe_0;
  wire  _T_1 = ~io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 72:17]
  assign mem_io_rdData_MPORT_en = mem_io_rdData_MPORT_en_pipe_0;
  assign mem_io_rdData_MPORT_addr = mem_io_rdData_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_io_rdData_MPORT_data = mem[mem_io_rdData_MPORT_addr]; // @[\\src\\main\\scala\\bram\\bramMem.scala 43:24]
  `else
  assign mem_io_rdData_MPORT_data = mem_io_rdData_MPORT_addr >= 5'h1c ? _RAND_1[27:0] : mem[mem_io_rdData_MPORT_addr]; // @[\\src\\main\\scala\\bram\\bramMem.scala 43:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = io_wrData;
  assign mem_MPORT_addr = io_addr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_en & io_wrEn;
  assign io_rdData = io_en & ~io_wrEn ? mem_io_rdData_MPORT_data : 28'h0; // @[\\src\\main\\scala\\bram\\bramMem.scala 71:13 72:27 73:13]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[\\src\\main\\scala\\bram\\bramMem.scala 43:24]
    end
    mem_io_rdData_MPORT_en_pipe_0 <= io_en & _T_1;
    if (io_en & _T_1) begin
      mem_io_rdData_MPORT_addr_pipe_0 <= io_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 28; initvar = initvar+1)
    mem[initvar] = _RAND_0[27:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_io_rdData_MPORT_en_pipe_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  mem_io_rdData_MPORT_addr_pipe_0 = _RAND_3[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BramMemWrapper(
  input         clock,
  input  [4:0]  io_lineAddr, // @[\\src\\main\\scala\\bram\\bramMem.scala 97:12]
  input         io_lineEn, // @[\\src\\main\\scala\\bram\\bramMem.scala 97:12]
  output [27:0] io_lineData, // @[\\src\\main\\scala\\bram\\bramMem.scala 97:12]
  input         io_wrEn, // @[\\src\\main\\scala\\bram\\bramMem.scala 97:12]
  input  [4:0]  io_wrAddr, // @[\\src\\main\\scala\\bram\\bramMem.scala 97:12]
  input  [27:0] io_wrData // @[\\src\\main\\scala\\bram\\bramMem.scala 97:12]
);
  wire  bramCore_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 110:22]
  wire [4:0] bramCore_io_addr; // @[\\src\\main\\scala\\bram\\bramMem.scala 110:22]
  wire  bramCore_io_en; // @[\\src\\main\\scala\\bram\\bramMem.scala 110:22]
  wire  bramCore_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 110:22]
  wire [27:0] bramCore_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 110:22]
  wire [27:0] bramCore_io_rdData; // @[\\src\\main\\scala\\bram\\bramMem.scala 110:22]
  BramMem bramCore ( // @[\\src\\main\\scala\\bram\\bramMem.scala 110:22]
    .clock(bramCore_clock),
    .io_addr(bramCore_io_addr),
    .io_en(bramCore_io_en),
    .io_wrEn(bramCore_io_wrEn),
    .io_wrData(bramCore_io_wrData),
    .io_rdData(bramCore_io_rdData)
  );
  assign io_lineData = bramCore_io_rdData; // @[\\src\\main\\scala\\bram\\bramMem.scala 122:13]
  assign bramCore_clock = clock;
  assign bramCore_io_addr = io_wrEn ? io_wrAddr : io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 118:24]
  assign bramCore_io_en = io_lineEn | io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 119:31]
  assign bramCore_io_wrEn = io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 113:20]
  assign bramCore_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 114:20]
endmodule
module t28x100(
  input         clock,
  input         reset,
  input  [4:0]  io_lineAddr, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  input         io_lineEn, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_0, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_1, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_2, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_3, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_4, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_5, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_6, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_7, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_8, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_9, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_10, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_11, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_12, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_13, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_14, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_15, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_16, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_17, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_18, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_19, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_20, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_21, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_22, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_23, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_24, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_25, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_26, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_27, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_28, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_29, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_30, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_31, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_32, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_33, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_34, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_35, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_36, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_37, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_38, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_39, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_40, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_41, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_42, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_43, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_44, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_45, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_46, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_47, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_48, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_49, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_50, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_51, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_52, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_53, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_54, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_55, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_56, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_57, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_58, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_59, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_60, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_61, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_62, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_63, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_64, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_65, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_66, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_67, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_68, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_69, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_70, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_71, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_72, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_73, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_74, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_75, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_76, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_77, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_78, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_79, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_80, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_81, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_82, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_83, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_84, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_85, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_86, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_87, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_88, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_89, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_90, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_91, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_92, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_93, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_94, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_95, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_96, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_97, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_98, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  output [27:0] io_lineData_99, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  input         io_wrEn, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  input  [6:0]  io_wrTemplate, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  input  [4:0]  io_wrAddr, // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
  input  [27:0] io_wrData // @[\\src\\main\\scala\\bram\\bramMem.scala 145:14]
);
  wire  templates_0_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_0_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_0_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_0_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_0_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_0_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_0_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_1_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_1_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_1_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_1_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_1_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_1_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_1_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_2_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_2_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_2_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_2_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_2_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_2_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_2_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_3_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_3_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_3_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_3_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_3_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_3_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_3_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_4_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_4_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_4_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_4_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_4_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_4_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_4_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_5_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_5_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_5_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_5_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_5_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_5_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_5_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_6_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_6_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_6_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_6_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_6_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_6_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_6_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_7_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_7_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_7_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_7_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_7_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_7_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_7_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_8_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_8_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_8_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_8_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_8_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_8_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_8_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_9_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_9_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_9_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_9_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_9_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_9_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_9_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_10_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_10_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_10_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_10_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_10_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_10_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_10_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_11_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_11_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_11_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_11_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_11_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_11_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_11_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_12_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_12_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_12_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_12_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_12_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_12_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_12_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_13_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_13_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_13_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_13_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_13_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_13_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_13_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_14_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_14_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_14_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_14_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_14_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_14_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_14_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_15_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_15_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_15_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_15_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_15_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_15_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_15_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_16_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_16_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_16_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_16_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_16_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_16_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_16_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_17_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_17_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_17_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_17_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_17_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_17_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_17_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_18_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_18_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_18_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_18_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_18_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_18_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_18_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_19_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_19_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_19_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_19_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_19_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_19_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_19_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_20_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_20_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_20_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_20_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_20_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_20_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_20_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_21_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_21_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_21_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_21_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_21_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_21_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_21_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_22_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_22_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_22_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_22_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_22_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_22_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_22_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_23_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_23_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_23_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_23_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_23_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_23_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_23_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_24_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_24_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_24_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_24_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_24_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_24_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_24_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_25_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_25_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_25_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_25_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_25_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_25_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_25_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_26_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_26_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_26_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_26_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_26_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_26_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_26_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_27_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_27_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_27_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_27_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_27_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_27_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_27_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_28_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_28_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_28_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_28_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_28_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_28_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_28_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_29_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_29_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_29_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_29_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_29_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_29_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_29_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_30_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_30_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_30_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_30_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_30_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_30_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_30_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_31_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_31_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_31_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_31_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_31_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_31_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_31_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_32_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_32_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_32_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_32_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_32_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_32_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_32_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_33_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_33_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_33_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_33_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_33_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_33_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_33_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_34_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_34_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_34_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_34_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_34_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_34_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_34_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_35_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_35_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_35_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_35_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_35_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_35_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_35_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_36_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_36_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_36_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_36_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_36_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_36_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_36_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_37_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_37_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_37_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_37_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_37_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_37_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_37_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_38_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_38_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_38_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_38_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_38_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_38_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_38_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_39_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_39_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_39_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_39_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_39_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_39_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_39_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_40_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_40_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_40_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_40_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_40_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_40_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_40_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_41_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_41_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_41_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_41_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_41_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_41_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_41_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_42_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_42_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_42_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_42_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_42_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_42_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_42_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_43_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_43_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_43_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_43_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_43_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_43_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_43_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_44_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_44_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_44_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_44_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_44_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_44_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_44_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_45_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_45_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_45_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_45_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_45_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_45_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_45_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_46_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_46_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_46_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_46_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_46_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_46_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_46_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_47_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_47_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_47_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_47_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_47_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_47_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_47_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_48_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_48_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_48_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_48_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_48_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_48_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_48_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_49_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_49_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_49_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_49_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_49_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_49_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_49_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_50_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_50_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_50_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_50_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_50_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_50_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_50_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_51_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_51_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_51_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_51_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_51_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_51_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_51_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_52_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_52_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_52_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_52_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_52_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_52_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_52_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_53_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_53_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_53_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_53_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_53_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_53_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_53_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_54_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_54_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_54_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_54_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_54_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_54_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_54_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_55_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_55_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_55_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_55_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_55_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_55_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_55_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_56_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_56_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_56_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_56_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_56_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_56_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_56_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_57_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_57_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_57_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_57_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_57_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_57_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_57_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_58_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_58_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_58_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_58_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_58_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_58_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_58_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_59_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_59_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_59_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_59_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_59_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_59_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_59_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_60_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_60_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_60_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_60_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_60_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_60_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_60_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_61_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_61_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_61_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_61_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_61_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_61_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_61_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_62_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_62_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_62_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_62_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_62_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_62_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_62_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_63_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_63_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_63_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_63_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_63_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_63_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_63_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_64_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_64_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_64_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_64_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_64_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_64_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_64_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_65_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_65_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_65_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_65_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_65_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_65_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_65_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_66_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_66_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_66_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_66_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_66_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_66_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_66_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_67_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_67_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_67_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_67_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_67_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_67_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_67_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_68_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_68_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_68_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_68_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_68_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_68_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_68_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_69_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_69_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_69_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_69_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_69_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_69_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_69_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_70_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_70_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_70_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_70_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_70_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_70_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_70_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_71_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_71_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_71_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_71_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_71_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_71_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_71_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_72_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_72_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_72_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_72_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_72_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_72_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_72_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_73_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_73_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_73_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_73_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_73_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_73_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_73_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_74_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_74_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_74_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_74_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_74_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_74_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_74_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_75_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_75_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_75_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_75_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_75_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_75_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_75_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_76_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_76_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_76_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_76_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_76_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_76_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_76_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_77_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_77_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_77_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_77_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_77_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_77_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_77_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_78_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_78_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_78_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_78_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_78_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_78_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_78_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_79_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_79_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_79_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_79_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_79_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_79_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_79_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_80_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_80_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_80_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_80_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_80_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_80_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_80_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_81_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_81_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_81_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_81_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_81_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_81_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_81_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_82_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_82_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_82_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_82_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_82_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_82_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_82_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_83_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_83_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_83_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_83_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_83_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_83_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_83_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_84_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_84_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_84_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_84_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_84_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_84_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_84_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_85_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_85_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_85_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_85_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_85_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_85_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_85_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_86_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_86_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_86_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_86_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_86_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_86_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_86_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_87_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_87_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_87_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_87_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_87_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_87_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_87_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_88_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_88_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_88_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_88_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_88_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_88_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_88_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_89_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_89_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_89_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_89_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_89_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_89_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_89_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_90_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_90_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_90_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_90_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_90_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_90_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_90_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_91_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_91_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_91_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_91_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_91_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_91_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_91_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_92_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_92_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_92_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_92_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_92_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_92_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_92_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_93_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_93_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_93_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_93_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_93_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_93_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_93_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_94_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_94_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_94_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_94_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_94_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_94_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_94_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_95_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_95_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_95_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_95_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_95_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_95_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_95_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_96_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_96_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_96_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_96_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_96_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_96_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_96_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_97_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_97_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_97_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_97_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_97_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_97_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_97_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_98_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_98_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_98_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_98_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_98_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_98_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_98_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_99_clock; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_99_io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_99_io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_99_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire  templates_99_io_wrEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [4:0] templates_99_io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  wire [27:0] templates_99_io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
  BramMemWrapper templates_0 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_0_clock),
    .io_lineAddr(templates_0_io_lineAddr),
    .io_lineEn(templates_0_io_lineEn),
    .io_lineData(templates_0_io_lineData),
    .io_wrEn(templates_0_io_wrEn),
    .io_wrAddr(templates_0_io_wrAddr),
    .io_wrData(templates_0_io_wrData)
  );
  BramMemWrapper templates_1 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_1_clock),
    .io_lineAddr(templates_1_io_lineAddr),
    .io_lineEn(templates_1_io_lineEn),
    .io_lineData(templates_1_io_lineData),
    .io_wrEn(templates_1_io_wrEn),
    .io_wrAddr(templates_1_io_wrAddr),
    .io_wrData(templates_1_io_wrData)
  );
  BramMemWrapper templates_2 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_2_clock),
    .io_lineAddr(templates_2_io_lineAddr),
    .io_lineEn(templates_2_io_lineEn),
    .io_lineData(templates_2_io_lineData),
    .io_wrEn(templates_2_io_wrEn),
    .io_wrAddr(templates_2_io_wrAddr),
    .io_wrData(templates_2_io_wrData)
  );
  BramMemWrapper templates_3 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_3_clock),
    .io_lineAddr(templates_3_io_lineAddr),
    .io_lineEn(templates_3_io_lineEn),
    .io_lineData(templates_3_io_lineData),
    .io_wrEn(templates_3_io_wrEn),
    .io_wrAddr(templates_3_io_wrAddr),
    .io_wrData(templates_3_io_wrData)
  );
  BramMemWrapper templates_4 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_4_clock),
    .io_lineAddr(templates_4_io_lineAddr),
    .io_lineEn(templates_4_io_lineEn),
    .io_lineData(templates_4_io_lineData),
    .io_wrEn(templates_4_io_wrEn),
    .io_wrAddr(templates_4_io_wrAddr),
    .io_wrData(templates_4_io_wrData)
  );
  BramMemWrapper templates_5 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_5_clock),
    .io_lineAddr(templates_5_io_lineAddr),
    .io_lineEn(templates_5_io_lineEn),
    .io_lineData(templates_5_io_lineData),
    .io_wrEn(templates_5_io_wrEn),
    .io_wrAddr(templates_5_io_wrAddr),
    .io_wrData(templates_5_io_wrData)
  );
  BramMemWrapper templates_6 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_6_clock),
    .io_lineAddr(templates_6_io_lineAddr),
    .io_lineEn(templates_6_io_lineEn),
    .io_lineData(templates_6_io_lineData),
    .io_wrEn(templates_6_io_wrEn),
    .io_wrAddr(templates_6_io_wrAddr),
    .io_wrData(templates_6_io_wrData)
  );
  BramMemWrapper templates_7 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_7_clock),
    .io_lineAddr(templates_7_io_lineAddr),
    .io_lineEn(templates_7_io_lineEn),
    .io_lineData(templates_7_io_lineData),
    .io_wrEn(templates_7_io_wrEn),
    .io_wrAddr(templates_7_io_wrAddr),
    .io_wrData(templates_7_io_wrData)
  );
  BramMemWrapper templates_8 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_8_clock),
    .io_lineAddr(templates_8_io_lineAddr),
    .io_lineEn(templates_8_io_lineEn),
    .io_lineData(templates_8_io_lineData),
    .io_wrEn(templates_8_io_wrEn),
    .io_wrAddr(templates_8_io_wrAddr),
    .io_wrData(templates_8_io_wrData)
  );
  BramMemWrapper templates_9 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_9_clock),
    .io_lineAddr(templates_9_io_lineAddr),
    .io_lineEn(templates_9_io_lineEn),
    .io_lineData(templates_9_io_lineData),
    .io_wrEn(templates_9_io_wrEn),
    .io_wrAddr(templates_9_io_wrAddr),
    .io_wrData(templates_9_io_wrData)
  );
  BramMemWrapper templates_10 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_10_clock),
    .io_lineAddr(templates_10_io_lineAddr),
    .io_lineEn(templates_10_io_lineEn),
    .io_lineData(templates_10_io_lineData),
    .io_wrEn(templates_10_io_wrEn),
    .io_wrAddr(templates_10_io_wrAddr),
    .io_wrData(templates_10_io_wrData)
  );
  BramMemWrapper templates_11 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_11_clock),
    .io_lineAddr(templates_11_io_lineAddr),
    .io_lineEn(templates_11_io_lineEn),
    .io_lineData(templates_11_io_lineData),
    .io_wrEn(templates_11_io_wrEn),
    .io_wrAddr(templates_11_io_wrAddr),
    .io_wrData(templates_11_io_wrData)
  );
  BramMemWrapper templates_12 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_12_clock),
    .io_lineAddr(templates_12_io_lineAddr),
    .io_lineEn(templates_12_io_lineEn),
    .io_lineData(templates_12_io_lineData),
    .io_wrEn(templates_12_io_wrEn),
    .io_wrAddr(templates_12_io_wrAddr),
    .io_wrData(templates_12_io_wrData)
  );
  BramMemWrapper templates_13 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_13_clock),
    .io_lineAddr(templates_13_io_lineAddr),
    .io_lineEn(templates_13_io_lineEn),
    .io_lineData(templates_13_io_lineData),
    .io_wrEn(templates_13_io_wrEn),
    .io_wrAddr(templates_13_io_wrAddr),
    .io_wrData(templates_13_io_wrData)
  );
  BramMemWrapper templates_14 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_14_clock),
    .io_lineAddr(templates_14_io_lineAddr),
    .io_lineEn(templates_14_io_lineEn),
    .io_lineData(templates_14_io_lineData),
    .io_wrEn(templates_14_io_wrEn),
    .io_wrAddr(templates_14_io_wrAddr),
    .io_wrData(templates_14_io_wrData)
  );
  BramMemWrapper templates_15 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_15_clock),
    .io_lineAddr(templates_15_io_lineAddr),
    .io_lineEn(templates_15_io_lineEn),
    .io_lineData(templates_15_io_lineData),
    .io_wrEn(templates_15_io_wrEn),
    .io_wrAddr(templates_15_io_wrAddr),
    .io_wrData(templates_15_io_wrData)
  );
  BramMemWrapper templates_16 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_16_clock),
    .io_lineAddr(templates_16_io_lineAddr),
    .io_lineEn(templates_16_io_lineEn),
    .io_lineData(templates_16_io_lineData),
    .io_wrEn(templates_16_io_wrEn),
    .io_wrAddr(templates_16_io_wrAddr),
    .io_wrData(templates_16_io_wrData)
  );
  BramMemWrapper templates_17 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_17_clock),
    .io_lineAddr(templates_17_io_lineAddr),
    .io_lineEn(templates_17_io_lineEn),
    .io_lineData(templates_17_io_lineData),
    .io_wrEn(templates_17_io_wrEn),
    .io_wrAddr(templates_17_io_wrAddr),
    .io_wrData(templates_17_io_wrData)
  );
  BramMemWrapper templates_18 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_18_clock),
    .io_lineAddr(templates_18_io_lineAddr),
    .io_lineEn(templates_18_io_lineEn),
    .io_lineData(templates_18_io_lineData),
    .io_wrEn(templates_18_io_wrEn),
    .io_wrAddr(templates_18_io_wrAddr),
    .io_wrData(templates_18_io_wrData)
  );
  BramMemWrapper templates_19 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_19_clock),
    .io_lineAddr(templates_19_io_lineAddr),
    .io_lineEn(templates_19_io_lineEn),
    .io_lineData(templates_19_io_lineData),
    .io_wrEn(templates_19_io_wrEn),
    .io_wrAddr(templates_19_io_wrAddr),
    .io_wrData(templates_19_io_wrData)
  );
  BramMemWrapper templates_20 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_20_clock),
    .io_lineAddr(templates_20_io_lineAddr),
    .io_lineEn(templates_20_io_lineEn),
    .io_lineData(templates_20_io_lineData),
    .io_wrEn(templates_20_io_wrEn),
    .io_wrAddr(templates_20_io_wrAddr),
    .io_wrData(templates_20_io_wrData)
  );
  BramMemWrapper templates_21 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_21_clock),
    .io_lineAddr(templates_21_io_lineAddr),
    .io_lineEn(templates_21_io_lineEn),
    .io_lineData(templates_21_io_lineData),
    .io_wrEn(templates_21_io_wrEn),
    .io_wrAddr(templates_21_io_wrAddr),
    .io_wrData(templates_21_io_wrData)
  );
  BramMemWrapper templates_22 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_22_clock),
    .io_lineAddr(templates_22_io_lineAddr),
    .io_lineEn(templates_22_io_lineEn),
    .io_lineData(templates_22_io_lineData),
    .io_wrEn(templates_22_io_wrEn),
    .io_wrAddr(templates_22_io_wrAddr),
    .io_wrData(templates_22_io_wrData)
  );
  BramMemWrapper templates_23 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_23_clock),
    .io_lineAddr(templates_23_io_lineAddr),
    .io_lineEn(templates_23_io_lineEn),
    .io_lineData(templates_23_io_lineData),
    .io_wrEn(templates_23_io_wrEn),
    .io_wrAddr(templates_23_io_wrAddr),
    .io_wrData(templates_23_io_wrData)
  );
  BramMemWrapper templates_24 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_24_clock),
    .io_lineAddr(templates_24_io_lineAddr),
    .io_lineEn(templates_24_io_lineEn),
    .io_lineData(templates_24_io_lineData),
    .io_wrEn(templates_24_io_wrEn),
    .io_wrAddr(templates_24_io_wrAddr),
    .io_wrData(templates_24_io_wrData)
  );
  BramMemWrapper templates_25 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_25_clock),
    .io_lineAddr(templates_25_io_lineAddr),
    .io_lineEn(templates_25_io_lineEn),
    .io_lineData(templates_25_io_lineData),
    .io_wrEn(templates_25_io_wrEn),
    .io_wrAddr(templates_25_io_wrAddr),
    .io_wrData(templates_25_io_wrData)
  );
  BramMemWrapper templates_26 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_26_clock),
    .io_lineAddr(templates_26_io_lineAddr),
    .io_lineEn(templates_26_io_lineEn),
    .io_lineData(templates_26_io_lineData),
    .io_wrEn(templates_26_io_wrEn),
    .io_wrAddr(templates_26_io_wrAddr),
    .io_wrData(templates_26_io_wrData)
  );
  BramMemWrapper templates_27 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_27_clock),
    .io_lineAddr(templates_27_io_lineAddr),
    .io_lineEn(templates_27_io_lineEn),
    .io_lineData(templates_27_io_lineData),
    .io_wrEn(templates_27_io_wrEn),
    .io_wrAddr(templates_27_io_wrAddr),
    .io_wrData(templates_27_io_wrData)
  );
  BramMemWrapper templates_28 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_28_clock),
    .io_lineAddr(templates_28_io_lineAddr),
    .io_lineEn(templates_28_io_lineEn),
    .io_lineData(templates_28_io_lineData),
    .io_wrEn(templates_28_io_wrEn),
    .io_wrAddr(templates_28_io_wrAddr),
    .io_wrData(templates_28_io_wrData)
  );
  BramMemWrapper templates_29 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_29_clock),
    .io_lineAddr(templates_29_io_lineAddr),
    .io_lineEn(templates_29_io_lineEn),
    .io_lineData(templates_29_io_lineData),
    .io_wrEn(templates_29_io_wrEn),
    .io_wrAddr(templates_29_io_wrAddr),
    .io_wrData(templates_29_io_wrData)
  );
  BramMemWrapper templates_30 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_30_clock),
    .io_lineAddr(templates_30_io_lineAddr),
    .io_lineEn(templates_30_io_lineEn),
    .io_lineData(templates_30_io_lineData),
    .io_wrEn(templates_30_io_wrEn),
    .io_wrAddr(templates_30_io_wrAddr),
    .io_wrData(templates_30_io_wrData)
  );
  BramMemWrapper templates_31 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_31_clock),
    .io_lineAddr(templates_31_io_lineAddr),
    .io_lineEn(templates_31_io_lineEn),
    .io_lineData(templates_31_io_lineData),
    .io_wrEn(templates_31_io_wrEn),
    .io_wrAddr(templates_31_io_wrAddr),
    .io_wrData(templates_31_io_wrData)
  );
  BramMemWrapper templates_32 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_32_clock),
    .io_lineAddr(templates_32_io_lineAddr),
    .io_lineEn(templates_32_io_lineEn),
    .io_lineData(templates_32_io_lineData),
    .io_wrEn(templates_32_io_wrEn),
    .io_wrAddr(templates_32_io_wrAddr),
    .io_wrData(templates_32_io_wrData)
  );
  BramMemWrapper templates_33 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_33_clock),
    .io_lineAddr(templates_33_io_lineAddr),
    .io_lineEn(templates_33_io_lineEn),
    .io_lineData(templates_33_io_lineData),
    .io_wrEn(templates_33_io_wrEn),
    .io_wrAddr(templates_33_io_wrAddr),
    .io_wrData(templates_33_io_wrData)
  );
  BramMemWrapper templates_34 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_34_clock),
    .io_lineAddr(templates_34_io_lineAddr),
    .io_lineEn(templates_34_io_lineEn),
    .io_lineData(templates_34_io_lineData),
    .io_wrEn(templates_34_io_wrEn),
    .io_wrAddr(templates_34_io_wrAddr),
    .io_wrData(templates_34_io_wrData)
  );
  BramMemWrapper templates_35 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_35_clock),
    .io_lineAddr(templates_35_io_lineAddr),
    .io_lineEn(templates_35_io_lineEn),
    .io_lineData(templates_35_io_lineData),
    .io_wrEn(templates_35_io_wrEn),
    .io_wrAddr(templates_35_io_wrAddr),
    .io_wrData(templates_35_io_wrData)
  );
  BramMemWrapper templates_36 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_36_clock),
    .io_lineAddr(templates_36_io_lineAddr),
    .io_lineEn(templates_36_io_lineEn),
    .io_lineData(templates_36_io_lineData),
    .io_wrEn(templates_36_io_wrEn),
    .io_wrAddr(templates_36_io_wrAddr),
    .io_wrData(templates_36_io_wrData)
  );
  BramMemWrapper templates_37 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_37_clock),
    .io_lineAddr(templates_37_io_lineAddr),
    .io_lineEn(templates_37_io_lineEn),
    .io_lineData(templates_37_io_lineData),
    .io_wrEn(templates_37_io_wrEn),
    .io_wrAddr(templates_37_io_wrAddr),
    .io_wrData(templates_37_io_wrData)
  );
  BramMemWrapper templates_38 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_38_clock),
    .io_lineAddr(templates_38_io_lineAddr),
    .io_lineEn(templates_38_io_lineEn),
    .io_lineData(templates_38_io_lineData),
    .io_wrEn(templates_38_io_wrEn),
    .io_wrAddr(templates_38_io_wrAddr),
    .io_wrData(templates_38_io_wrData)
  );
  BramMemWrapper templates_39 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_39_clock),
    .io_lineAddr(templates_39_io_lineAddr),
    .io_lineEn(templates_39_io_lineEn),
    .io_lineData(templates_39_io_lineData),
    .io_wrEn(templates_39_io_wrEn),
    .io_wrAddr(templates_39_io_wrAddr),
    .io_wrData(templates_39_io_wrData)
  );
  BramMemWrapper templates_40 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_40_clock),
    .io_lineAddr(templates_40_io_lineAddr),
    .io_lineEn(templates_40_io_lineEn),
    .io_lineData(templates_40_io_lineData),
    .io_wrEn(templates_40_io_wrEn),
    .io_wrAddr(templates_40_io_wrAddr),
    .io_wrData(templates_40_io_wrData)
  );
  BramMemWrapper templates_41 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_41_clock),
    .io_lineAddr(templates_41_io_lineAddr),
    .io_lineEn(templates_41_io_lineEn),
    .io_lineData(templates_41_io_lineData),
    .io_wrEn(templates_41_io_wrEn),
    .io_wrAddr(templates_41_io_wrAddr),
    .io_wrData(templates_41_io_wrData)
  );
  BramMemWrapper templates_42 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_42_clock),
    .io_lineAddr(templates_42_io_lineAddr),
    .io_lineEn(templates_42_io_lineEn),
    .io_lineData(templates_42_io_lineData),
    .io_wrEn(templates_42_io_wrEn),
    .io_wrAddr(templates_42_io_wrAddr),
    .io_wrData(templates_42_io_wrData)
  );
  BramMemWrapper templates_43 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_43_clock),
    .io_lineAddr(templates_43_io_lineAddr),
    .io_lineEn(templates_43_io_lineEn),
    .io_lineData(templates_43_io_lineData),
    .io_wrEn(templates_43_io_wrEn),
    .io_wrAddr(templates_43_io_wrAddr),
    .io_wrData(templates_43_io_wrData)
  );
  BramMemWrapper templates_44 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_44_clock),
    .io_lineAddr(templates_44_io_lineAddr),
    .io_lineEn(templates_44_io_lineEn),
    .io_lineData(templates_44_io_lineData),
    .io_wrEn(templates_44_io_wrEn),
    .io_wrAddr(templates_44_io_wrAddr),
    .io_wrData(templates_44_io_wrData)
  );
  BramMemWrapper templates_45 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_45_clock),
    .io_lineAddr(templates_45_io_lineAddr),
    .io_lineEn(templates_45_io_lineEn),
    .io_lineData(templates_45_io_lineData),
    .io_wrEn(templates_45_io_wrEn),
    .io_wrAddr(templates_45_io_wrAddr),
    .io_wrData(templates_45_io_wrData)
  );
  BramMemWrapper templates_46 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_46_clock),
    .io_lineAddr(templates_46_io_lineAddr),
    .io_lineEn(templates_46_io_lineEn),
    .io_lineData(templates_46_io_lineData),
    .io_wrEn(templates_46_io_wrEn),
    .io_wrAddr(templates_46_io_wrAddr),
    .io_wrData(templates_46_io_wrData)
  );
  BramMemWrapper templates_47 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_47_clock),
    .io_lineAddr(templates_47_io_lineAddr),
    .io_lineEn(templates_47_io_lineEn),
    .io_lineData(templates_47_io_lineData),
    .io_wrEn(templates_47_io_wrEn),
    .io_wrAddr(templates_47_io_wrAddr),
    .io_wrData(templates_47_io_wrData)
  );
  BramMemWrapper templates_48 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_48_clock),
    .io_lineAddr(templates_48_io_lineAddr),
    .io_lineEn(templates_48_io_lineEn),
    .io_lineData(templates_48_io_lineData),
    .io_wrEn(templates_48_io_wrEn),
    .io_wrAddr(templates_48_io_wrAddr),
    .io_wrData(templates_48_io_wrData)
  );
  BramMemWrapper templates_49 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_49_clock),
    .io_lineAddr(templates_49_io_lineAddr),
    .io_lineEn(templates_49_io_lineEn),
    .io_lineData(templates_49_io_lineData),
    .io_wrEn(templates_49_io_wrEn),
    .io_wrAddr(templates_49_io_wrAddr),
    .io_wrData(templates_49_io_wrData)
  );
  BramMemWrapper templates_50 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_50_clock),
    .io_lineAddr(templates_50_io_lineAddr),
    .io_lineEn(templates_50_io_lineEn),
    .io_lineData(templates_50_io_lineData),
    .io_wrEn(templates_50_io_wrEn),
    .io_wrAddr(templates_50_io_wrAddr),
    .io_wrData(templates_50_io_wrData)
  );
  BramMemWrapper templates_51 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_51_clock),
    .io_lineAddr(templates_51_io_lineAddr),
    .io_lineEn(templates_51_io_lineEn),
    .io_lineData(templates_51_io_lineData),
    .io_wrEn(templates_51_io_wrEn),
    .io_wrAddr(templates_51_io_wrAddr),
    .io_wrData(templates_51_io_wrData)
  );
  BramMemWrapper templates_52 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_52_clock),
    .io_lineAddr(templates_52_io_lineAddr),
    .io_lineEn(templates_52_io_lineEn),
    .io_lineData(templates_52_io_lineData),
    .io_wrEn(templates_52_io_wrEn),
    .io_wrAddr(templates_52_io_wrAddr),
    .io_wrData(templates_52_io_wrData)
  );
  BramMemWrapper templates_53 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_53_clock),
    .io_lineAddr(templates_53_io_lineAddr),
    .io_lineEn(templates_53_io_lineEn),
    .io_lineData(templates_53_io_lineData),
    .io_wrEn(templates_53_io_wrEn),
    .io_wrAddr(templates_53_io_wrAddr),
    .io_wrData(templates_53_io_wrData)
  );
  BramMemWrapper templates_54 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_54_clock),
    .io_lineAddr(templates_54_io_lineAddr),
    .io_lineEn(templates_54_io_lineEn),
    .io_lineData(templates_54_io_lineData),
    .io_wrEn(templates_54_io_wrEn),
    .io_wrAddr(templates_54_io_wrAddr),
    .io_wrData(templates_54_io_wrData)
  );
  BramMemWrapper templates_55 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_55_clock),
    .io_lineAddr(templates_55_io_lineAddr),
    .io_lineEn(templates_55_io_lineEn),
    .io_lineData(templates_55_io_lineData),
    .io_wrEn(templates_55_io_wrEn),
    .io_wrAddr(templates_55_io_wrAddr),
    .io_wrData(templates_55_io_wrData)
  );
  BramMemWrapper templates_56 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_56_clock),
    .io_lineAddr(templates_56_io_lineAddr),
    .io_lineEn(templates_56_io_lineEn),
    .io_lineData(templates_56_io_lineData),
    .io_wrEn(templates_56_io_wrEn),
    .io_wrAddr(templates_56_io_wrAddr),
    .io_wrData(templates_56_io_wrData)
  );
  BramMemWrapper templates_57 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_57_clock),
    .io_lineAddr(templates_57_io_lineAddr),
    .io_lineEn(templates_57_io_lineEn),
    .io_lineData(templates_57_io_lineData),
    .io_wrEn(templates_57_io_wrEn),
    .io_wrAddr(templates_57_io_wrAddr),
    .io_wrData(templates_57_io_wrData)
  );
  BramMemWrapper templates_58 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_58_clock),
    .io_lineAddr(templates_58_io_lineAddr),
    .io_lineEn(templates_58_io_lineEn),
    .io_lineData(templates_58_io_lineData),
    .io_wrEn(templates_58_io_wrEn),
    .io_wrAddr(templates_58_io_wrAddr),
    .io_wrData(templates_58_io_wrData)
  );
  BramMemWrapper templates_59 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_59_clock),
    .io_lineAddr(templates_59_io_lineAddr),
    .io_lineEn(templates_59_io_lineEn),
    .io_lineData(templates_59_io_lineData),
    .io_wrEn(templates_59_io_wrEn),
    .io_wrAddr(templates_59_io_wrAddr),
    .io_wrData(templates_59_io_wrData)
  );
  BramMemWrapper templates_60 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_60_clock),
    .io_lineAddr(templates_60_io_lineAddr),
    .io_lineEn(templates_60_io_lineEn),
    .io_lineData(templates_60_io_lineData),
    .io_wrEn(templates_60_io_wrEn),
    .io_wrAddr(templates_60_io_wrAddr),
    .io_wrData(templates_60_io_wrData)
  );
  BramMemWrapper templates_61 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_61_clock),
    .io_lineAddr(templates_61_io_lineAddr),
    .io_lineEn(templates_61_io_lineEn),
    .io_lineData(templates_61_io_lineData),
    .io_wrEn(templates_61_io_wrEn),
    .io_wrAddr(templates_61_io_wrAddr),
    .io_wrData(templates_61_io_wrData)
  );
  BramMemWrapper templates_62 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_62_clock),
    .io_lineAddr(templates_62_io_lineAddr),
    .io_lineEn(templates_62_io_lineEn),
    .io_lineData(templates_62_io_lineData),
    .io_wrEn(templates_62_io_wrEn),
    .io_wrAddr(templates_62_io_wrAddr),
    .io_wrData(templates_62_io_wrData)
  );
  BramMemWrapper templates_63 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_63_clock),
    .io_lineAddr(templates_63_io_lineAddr),
    .io_lineEn(templates_63_io_lineEn),
    .io_lineData(templates_63_io_lineData),
    .io_wrEn(templates_63_io_wrEn),
    .io_wrAddr(templates_63_io_wrAddr),
    .io_wrData(templates_63_io_wrData)
  );
  BramMemWrapper templates_64 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_64_clock),
    .io_lineAddr(templates_64_io_lineAddr),
    .io_lineEn(templates_64_io_lineEn),
    .io_lineData(templates_64_io_lineData),
    .io_wrEn(templates_64_io_wrEn),
    .io_wrAddr(templates_64_io_wrAddr),
    .io_wrData(templates_64_io_wrData)
  );
  BramMemWrapper templates_65 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_65_clock),
    .io_lineAddr(templates_65_io_lineAddr),
    .io_lineEn(templates_65_io_lineEn),
    .io_lineData(templates_65_io_lineData),
    .io_wrEn(templates_65_io_wrEn),
    .io_wrAddr(templates_65_io_wrAddr),
    .io_wrData(templates_65_io_wrData)
  );
  BramMemWrapper templates_66 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_66_clock),
    .io_lineAddr(templates_66_io_lineAddr),
    .io_lineEn(templates_66_io_lineEn),
    .io_lineData(templates_66_io_lineData),
    .io_wrEn(templates_66_io_wrEn),
    .io_wrAddr(templates_66_io_wrAddr),
    .io_wrData(templates_66_io_wrData)
  );
  BramMemWrapper templates_67 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_67_clock),
    .io_lineAddr(templates_67_io_lineAddr),
    .io_lineEn(templates_67_io_lineEn),
    .io_lineData(templates_67_io_lineData),
    .io_wrEn(templates_67_io_wrEn),
    .io_wrAddr(templates_67_io_wrAddr),
    .io_wrData(templates_67_io_wrData)
  );
  BramMemWrapper templates_68 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_68_clock),
    .io_lineAddr(templates_68_io_lineAddr),
    .io_lineEn(templates_68_io_lineEn),
    .io_lineData(templates_68_io_lineData),
    .io_wrEn(templates_68_io_wrEn),
    .io_wrAddr(templates_68_io_wrAddr),
    .io_wrData(templates_68_io_wrData)
  );
  BramMemWrapper templates_69 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_69_clock),
    .io_lineAddr(templates_69_io_lineAddr),
    .io_lineEn(templates_69_io_lineEn),
    .io_lineData(templates_69_io_lineData),
    .io_wrEn(templates_69_io_wrEn),
    .io_wrAddr(templates_69_io_wrAddr),
    .io_wrData(templates_69_io_wrData)
  );
  BramMemWrapper templates_70 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_70_clock),
    .io_lineAddr(templates_70_io_lineAddr),
    .io_lineEn(templates_70_io_lineEn),
    .io_lineData(templates_70_io_lineData),
    .io_wrEn(templates_70_io_wrEn),
    .io_wrAddr(templates_70_io_wrAddr),
    .io_wrData(templates_70_io_wrData)
  );
  BramMemWrapper templates_71 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_71_clock),
    .io_lineAddr(templates_71_io_lineAddr),
    .io_lineEn(templates_71_io_lineEn),
    .io_lineData(templates_71_io_lineData),
    .io_wrEn(templates_71_io_wrEn),
    .io_wrAddr(templates_71_io_wrAddr),
    .io_wrData(templates_71_io_wrData)
  );
  BramMemWrapper templates_72 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_72_clock),
    .io_lineAddr(templates_72_io_lineAddr),
    .io_lineEn(templates_72_io_lineEn),
    .io_lineData(templates_72_io_lineData),
    .io_wrEn(templates_72_io_wrEn),
    .io_wrAddr(templates_72_io_wrAddr),
    .io_wrData(templates_72_io_wrData)
  );
  BramMemWrapper templates_73 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_73_clock),
    .io_lineAddr(templates_73_io_lineAddr),
    .io_lineEn(templates_73_io_lineEn),
    .io_lineData(templates_73_io_lineData),
    .io_wrEn(templates_73_io_wrEn),
    .io_wrAddr(templates_73_io_wrAddr),
    .io_wrData(templates_73_io_wrData)
  );
  BramMemWrapper templates_74 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_74_clock),
    .io_lineAddr(templates_74_io_lineAddr),
    .io_lineEn(templates_74_io_lineEn),
    .io_lineData(templates_74_io_lineData),
    .io_wrEn(templates_74_io_wrEn),
    .io_wrAddr(templates_74_io_wrAddr),
    .io_wrData(templates_74_io_wrData)
  );
  BramMemWrapper templates_75 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_75_clock),
    .io_lineAddr(templates_75_io_lineAddr),
    .io_lineEn(templates_75_io_lineEn),
    .io_lineData(templates_75_io_lineData),
    .io_wrEn(templates_75_io_wrEn),
    .io_wrAddr(templates_75_io_wrAddr),
    .io_wrData(templates_75_io_wrData)
  );
  BramMemWrapper templates_76 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_76_clock),
    .io_lineAddr(templates_76_io_lineAddr),
    .io_lineEn(templates_76_io_lineEn),
    .io_lineData(templates_76_io_lineData),
    .io_wrEn(templates_76_io_wrEn),
    .io_wrAddr(templates_76_io_wrAddr),
    .io_wrData(templates_76_io_wrData)
  );
  BramMemWrapper templates_77 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_77_clock),
    .io_lineAddr(templates_77_io_lineAddr),
    .io_lineEn(templates_77_io_lineEn),
    .io_lineData(templates_77_io_lineData),
    .io_wrEn(templates_77_io_wrEn),
    .io_wrAddr(templates_77_io_wrAddr),
    .io_wrData(templates_77_io_wrData)
  );
  BramMemWrapper templates_78 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_78_clock),
    .io_lineAddr(templates_78_io_lineAddr),
    .io_lineEn(templates_78_io_lineEn),
    .io_lineData(templates_78_io_lineData),
    .io_wrEn(templates_78_io_wrEn),
    .io_wrAddr(templates_78_io_wrAddr),
    .io_wrData(templates_78_io_wrData)
  );
  BramMemWrapper templates_79 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_79_clock),
    .io_lineAddr(templates_79_io_lineAddr),
    .io_lineEn(templates_79_io_lineEn),
    .io_lineData(templates_79_io_lineData),
    .io_wrEn(templates_79_io_wrEn),
    .io_wrAddr(templates_79_io_wrAddr),
    .io_wrData(templates_79_io_wrData)
  );
  BramMemWrapper templates_80 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_80_clock),
    .io_lineAddr(templates_80_io_lineAddr),
    .io_lineEn(templates_80_io_lineEn),
    .io_lineData(templates_80_io_lineData),
    .io_wrEn(templates_80_io_wrEn),
    .io_wrAddr(templates_80_io_wrAddr),
    .io_wrData(templates_80_io_wrData)
  );
  BramMemWrapper templates_81 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_81_clock),
    .io_lineAddr(templates_81_io_lineAddr),
    .io_lineEn(templates_81_io_lineEn),
    .io_lineData(templates_81_io_lineData),
    .io_wrEn(templates_81_io_wrEn),
    .io_wrAddr(templates_81_io_wrAddr),
    .io_wrData(templates_81_io_wrData)
  );
  BramMemWrapper templates_82 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_82_clock),
    .io_lineAddr(templates_82_io_lineAddr),
    .io_lineEn(templates_82_io_lineEn),
    .io_lineData(templates_82_io_lineData),
    .io_wrEn(templates_82_io_wrEn),
    .io_wrAddr(templates_82_io_wrAddr),
    .io_wrData(templates_82_io_wrData)
  );
  BramMemWrapper templates_83 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_83_clock),
    .io_lineAddr(templates_83_io_lineAddr),
    .io_lineEn(templates_83_io_lineEn),
    .io_lineData(templates_83_io_lineData),
    .io_wrEn(templates_83_io_wrEn),
    .io_wrAddr(templates_83_io_wrAddr),
    .io_wrData(templates_83_io_wrData)
  );
  BramMemWrapper templates_84 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_84_clock),
    .io_lineAddr(templates_84_io_lineAddr),
    .io_lineEn(templates_84_io_lineEn),
    .io_lineData(templates_84_io_lineData),
    .io_wrEn(templates_84_io_wrEn),
    .io_wrAddr(templates_84_io_wrAddr),
    .io_wrData(templates_84_io_wrData)
  );
  BramMemWrapper templates_85 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_85_clock),
    .io_lineAddr(templates_85_io_lineAddr),
    .io_lineEn(templates_85_io_lineEn),
    .io_lineData(templates_85_io_lineData),
    .io_wrEn(templates_85_io_wrEn),
    .io_wrAddr(templates_85_io_wrAddr),
    .io_wrData(templates_85_io_wrData)
  );
  BramMemWrapper templates_86 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_86_clock),
    .io_lineAddr(templates_86_io_lineAddr),
    .io_lineEn(templates_86_io_lineEn),
    .io_lineData(templates_86_io_lineData),
    .io_wrEn(templates_86_io_wrEn),
    .io_wrAddr(templates_86_io_wrAddr),
    .io_wrData(templates_86_io_wrData)
  );
  BramMemWrapper templates_87 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_87_clock),
    .io_lineAddr(templates_87_io_lineAddr),
    .io_lineEn(templates_87_io_lineEn),
    .io_lineData(templates_87_io_lineData),
    .io_wrEn(templates_87_io_wrEn),
    .io_wrAddr(templates_87_io_wrAddr),
    .io_wrData(templates_87_io_wrData)
  );
  BramMemWrapper templates_88 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_88_clock),
    .io_lineAddr(templates_88_io_lineAddr),
    .io_lineEn(templates_88_io_lineEn),
    .io_lineData(templates_88_io_lineData),
    .io_wrEn(templates_88_io_wrEn),
    .io_wrAddr(templates_88_io_wrAddr),
    .io_wrData(templates_88_io_wrData)
  );
  BramMemWrapper templates_89 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_89_clock),
    .io_lineAddr(templates_89_io_lineAddr),
    .io_lineEn(templates_89_io_lineEn),
    .io_lineData(templates_89_io_lineData),
    .io_wrEn(templates_89_io_wrEn),
    .io_wrAddr(templates_89_io_wrAddr),
    .io_wrData(templates_89_io_wrData)
  );
  BramMemWrapper templates_90 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_90_clock),
    .io_lineAddr(templates_90_io_lineAddr),
    .io_lineEn(templates_90_io_lineEn),
    .io_lineData(templates_90_io_lineData),
    .io_wrEn(templates_90_io_wrEn),
    .io_wrAddr(templates_90_io_wrAddr),
    .io_wrData(templates_90_io_wrData)
  );
  BramMemWrapper templates_91 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_91_clock),
    .io_lineAddr(templates_91_io_lineAddr),
    .io_lineEn(templates_91_io_lineEn),
    .io_lineData(templates_91_io_lineData),
    .io_wrEn(templates_91_io_wrEn),
    .io_wrAddr(templates_91_io_wrAddr),
    .io_wrData(templates_91_io_wrData)
  );
  BramMemWrapper templates_92 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_92_clock),
    .io_lineAddr(templates_92_io_lineAddr),
    .io_lineEn(templates_92_io_lineEn),
    .io_lineData(templates_92_io_lineData),
    .io_wrEn(templates_92_io_wrEn),
    .io_wrAddr(templates_92_io_wrAddr),
    .io_wrData(templates_92_io_wrData)
  );
  BramMemWrapper templates_93 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_93_clock),
    .io_lineAddr(templates_93_io_lineAddr),
    .io_lineEn(templates_93_io_lineEn),
    .io_lineData(templates_93_io_lineData),
    .io_wrEn(templates_93_io_wrEn),
    .io_wrAddr(templates_93_io_wrAddr),
    .io_wrData(templates_93_io_wrData)
  );
  BramMemWrapper templates_94 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_94_clock),
    .io_lineAddr(templates_94_io_lineAddr),
    .io_lineEn(templates_94_io_lineEn),
    .io_lineData(templates_94_io_lineData),
    .io_wrEn(templates_94_io_wrEn),
    .io_wrAddr(templates_94_io_wrAddr),
    .io_wrData(templates_94_io_wrData)
  );
  BramMemWrapper templates_95 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_95_clock),
    .io_lineAddr(templates_95_io_lineAddr),
    .io_lineEn(templates_95_io_lineEn),
    .io_lineData(templates_95_io_lineData),
    .io_wrEn(templates_95_io_wrEn),
    .io_wrAddr(templates_95_io_wrAddr),
    .io_wrData(templates_95_io_wrData)
  );
  BramMemWrapper templates_96 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_96_clock),
    .io_lineAddr(templates_96_io_lineAddr),
    .io_lineEn(templates_96_io_lineEn),
    .io_lineData(templates_96_io_lineData),
    .io_wrEn(templates_96_io_wrEn),
    .io_wrAddr(templates_96_io_wrAddr),
    .io_wrData(templates_96_io_wrData)
  );
  BramMemWrapper templates_97 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_97_clock),
    .io_lineAddr(templates_97_io_lineAddr),
    .io_lineEn(templates_97_io_lineEn),
    .io_lineData(templates_97_io_lineData),
    .io_wrEn(templates_97_io_wrEn),
    .io_wrAddr(templates_97_io_wrAddr),
    .io_wrData(templates_97_io_wrData)
  );
  BramMemWrapper templates_98 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_98_clock),
    .io_lineAddr(templates_98_io_lineAddr),
    .io_lineEn(templates_98_io_lineEn),
    .io_lineData(templates_98_io_lineData),
    .io_wrEn(templates_98_io_wrEn),
    .io_wrAddr(templates_98_io_wrAddr),
    .io_wrData(templates_98_io_wrData)
  );
  BramMemWrapper templates_99 ( // @[\\src\\main\\scala\\bram\\bramMem.scala 172:36]
    .clock(templates_99_clock),
    .io_lineAddr(templates_99_io_lineAddr),
    .io_lineEn(templates_99_io_lineEn),
    .io_lineData(templates_99_io_lineData),
    .io_wrEn(templates_99_io_wrEn),
    .io_wrAddr(templates_99_io_wrAddr),
    .io_wrData(templates_99_io_wrData)
  );
  assign io_lineData_0 = templates_0_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_1 = templates_1_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_2 = templates_2_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_3 = templates_3_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_4 = templates_4_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_5 = templates_5_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_6 = templates_6_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_7 = templates_7_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_8 = templates_8_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_9 = templates_9_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_10 = templates_10_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_11 = templates_11_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_12 = templates_12_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_13 = templates_13_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_14 = templates_14_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_15 = templates_15_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_16 = templates_16_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_17 = templates_17_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_18 = templates_18_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_19 = templates_19_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_20 = templates_20_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_21 = templates_21_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_22 = templates_22_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_23 = templates_23_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_24 = templates_24_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_25 = templates_25_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_26 = templates_26_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_27 = templates_27_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_28 = templates_28_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_29 = templates_29_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_30 = templates_30_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_31 = templates_31_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_32 = templates_32_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_33 = templates_33_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_34 = templates_34_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_35 = templates_35_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_36 = templates_36_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_37 = templates_37_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_38 = templates_38_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_39 = templates_39_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_40 = templates_40_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_41 = templates_41_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_42 = templates_42_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_43 = templates_43_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_44 = templates_44_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_45 = templates_45_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_46 = templates_46_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_47 = templates_47_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_48 = templates_48_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_49 = templates_49_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_50 = templates_50_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_51 = templates_51_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_52 = templates_52_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_53 = templates_53_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_54 = templates_54_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_55 = templates_55_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_56 = templates_56_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_57 = templates_57_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_58 = templates_58_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_59 = templates_59_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_60 = templates_60_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_61 = templates_61_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_62 = templates_62_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_63 = templates_63_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_64 = templates_64_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_65 = templates_65_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_66 = templates_66_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_67 = templates_67_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_68 = templates_68_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_69 = templates_69_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_70 = templates_70_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_71 = templates_71_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_72 = templates_72_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_73 = templates_73_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_74 = templates_74_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_75 = templates_75_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_76 = templates_76_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_77 = templates_77_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_78 = templates_78_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_79 = templates_79_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_80 = templates_80_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_81 = templates_81_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_82 = templates_82_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_83 = templates_83_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_84 = templates_84_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_85 = templates_85_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_86 = templates_86_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_87 = templates_87_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_88 = templates_88_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_89 = templates_89_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_90 = templates_90_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_91 = templates_91_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_92 = templates_92_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_93 = templates_93_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_94 = templates_94_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_95 = templates_95_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_96 = templates_96_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_97 = templates_97_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_98 = templates_98_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign io_lineData_99 = templates_99_io_lineData; // @[\\src\\main\\scala\\bram\\bramMem.scala 180:34]
  assign templates_0_clock = clock;
  assign templates_0_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_0_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_0_io_wrEn = io_wrEn & io_wrTemplate == 7'h0; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_0_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_0_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_1_clock = clock;
  assign templates_1_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_1_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_1_io_wrEn = io_wrEn & io_wrTemplate == 7'h1; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_1_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_1_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_2_clock = clock;
  assign templates_2_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_2_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_2_io_wrEn = io_wrEn & io_wrTemplate == 7'h2; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_2_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_2_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_3_clock = clock;
  assign templates_3_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_3_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_3_io_wrEn = io_wrEn & io_wrTemplate == 7'h3; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_3_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_3_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_4_clock = clock;
  assign templates_4_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_4_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_4_io_wrEn = io_wrEn & io_wrTemplate == 7'h4; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_4_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_4_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_5_clock = clock;
  assign templates_5_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_5_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_5_io_wrEn = io_wrEn & io_wrTemplate == 7'h5; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_5_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_5_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_6_clock = clock;
  assign templates_6_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_6_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_6_io_wrEn = io_wrEn & io_wrTemplate == 7'h6; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_6_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_6_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_7_clock = clock;
  assign templates_7_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_7_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_7_io_wrEn = io_wrEn & io_wrTemplate == 7'h7; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_7_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_7_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_8_clock = clock;
  assign templates_8_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_8_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_8_io_wrEn = io_wrEn & io_wrTemplate == 7'h8; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_8_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_8_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_9_clock = clock;
  assign templates_9_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_9_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_9_io_wrEn = io_wrEn & io_wrTemplate == 7'h9; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_9_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_9_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_10_clock = clock;
  assign templates_10_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_10_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_10_io_wrEn = io_wrEn & io_wrTemplate == 7'ha; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_10_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_10_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_11_clock = clock;
  assign templates_11_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_11_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_11_io_wrEn = io_wrEn & io_wrTemplate == 7'hb; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_11_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_11_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_12_clock = clock;
  assign templates_12_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_12_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_12_io_wrEn = io_wrEn & io_wrTemplate == 7'hc; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_12_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_12_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_13_clock = clock;
  assign templates_13_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_13_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_13_io_wrEn = io_wrEn & io_wrTemplate == 7'hd; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_13_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_13_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_14_clock = clock;
  assign templates_14_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_14_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_14_io_wrEn = io_wrEn & io_wrTemplate == 7'he; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_14_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_14_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_15_clock = clock;
  assign templates_15_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_15_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_15_io_wrEn = io_wrEn & io_wrTemplate == 7'hf; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_15_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_15_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_16_clock = clock;
  assign templates_16_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_16_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_16_io_wrEn = io_wrEn & io_wrTemplate == 7'h10; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_16_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_16_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_17_clock = clock;
  assign templates_17_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_17_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_17_io_wrEn = io_wrEn & io_wrTemplate == 7'h11; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_17_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_17_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_18_clock = clock;
  assign templates_18_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_18_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_18_io_wrEn = io_wrEn & io_wrTemplate == 7'h12; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_18_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_18_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_19_clock = clock;
  assign templates_19_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_19_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_19_io_wrEn = io_wrEn & io_wrTemplate == 7'h13; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_19_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_19_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_20_clock = clock;
  assign templates_20_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_20_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_20_io_wrEn = io_wrEn & io_wrTemplate == 7'h14; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_20_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_20_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_21_clock = clock;
  assign templates_21_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_21_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_21_io_wrEn = io_wrEn & io_wrTemplate == 7'h15; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_21_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_21_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_22_clock = clock;
  assign templates_22_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_22_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_22_io_wrEn = io_wrEn & io_wrTemplate == 7'h16; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_22_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_22_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_23_clock = clock;
  assign templates_23_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_23_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_23_io_wrEn = io_wrEn & io_wrTemplate == 7'h17; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_23_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_23_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_24_clock = clock;
  assign templates_24_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_24_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_24_io_wrEn = io_wrEn & io_wrTemplate == 7'h18; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_24_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_24_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_25_clock = clock;
  assign templates_25_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_25_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_25_io_wrEn = io_wrEn & io_wrTemplate == 7'h19; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_25_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_25_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_26_clock = clock;
  assign templates_26_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_26_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_26_io_wrEn = io_wrEn & io_wrTemplate == 7'h1a; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_26_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_26_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_27_clock = clock;
  assign templates_27_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_27_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_27_io_wrEn = io_wrEn & io_wrTemplate == 7'h1b; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_27_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_27_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_28_clock = clock;
  assign templates_28_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_28_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_28_io_wrEn = io_wrEn & io_wrTemplate == 7'h1c; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_28_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_28_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_29_clock = clock;
  assign templates_29_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_29_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_29_io_wrEn = io_wrEn & io_wrTemplate == 7'h1d; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_29_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_29_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_30_clock = clock;
  assign templates_30_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_30_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_30_io_wrEn = io_wrEn & io_wrTemplate == 7'h1e; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_30_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_30_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_31_clock = clock;
  assign templates_31_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_31_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_31_io_wrEn = io_wrEn & io_wrTemplate == 7'h1f; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_31_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_31_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_32_clock = clock;
  assign templates_32_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_32_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_32_io_wrEn = io_wrEn & io_wrTemplate == 7'h20; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_32_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_32_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_33_clock = clock;
  assign templates_33_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_33_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_33_io_wrEn = io_wrEn & io_wrTemplate == 7'h21; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_33_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_33_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_34_clock = clock;
  assign templates_34_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_34_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_34_io_wrEn = io_wrEn & io_wrTemplate == 7'h22; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_34_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_34_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_35_clock = clock;
  assign templates_35_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_35_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_35_io_wrEn = io_wrEn & io_wrTemplate == 7'h23; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_35_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_35_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_36_clock = clock;
  assign templates_36_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_36_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_36_io_wrEn = io_wrEn & io_wrTemplate == 7'h24; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_36_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_36_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_37_clock = clock;
  assign templates_37_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_37_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_37_io_wrEn = io_wrEn & io_wrTemplate == 7'h25; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_37_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_37_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_38_clock = clock;
  assign templates_38_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_38_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_38_io_wrEn = io_wrEn & io_wrTemplate == 7'h26; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_38_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_38_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_39_clock = clock;
  assign templates_39_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_39_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_39_io_wrEn = io_wrEn & io_wrTemplate == 7'h27; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_39_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_39_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_40_clock = clock;
  assign templates_40_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_40_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_40_io_wrEn = io_wrEn & io_wrTemplate == 7'h28; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_40_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_40_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_41_clock = clock;
  assign templates_41_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_41_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_41_io_wrEn = io_wrEn & io_wrTemplate == 7'h29; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_41_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_41_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_42_clock = clock;
  assign templates_42_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_42_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_42_io_wrEn = io_wrEn & io_wrTemplate == 7'h2a; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_42_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_42_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_43_clock = clock;
  assign templates_43_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_43_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_43_io_wrEn = io_wrEn & io_wrTemplate == 7'h2b; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_43_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_43_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_44_clock = clock;
  assign templates_44_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_44_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_44_io_wrEn = io_wrEn & io_wrTemplate == 7'h2c; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_44_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_44_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_45_clock = clock;
  assign templates_45_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_45_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_45_io_wrEn = io_wrEn & io_wrTemplate == 7'h2d; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_45_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_45_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_46_clock = clock;
  assign templates_46_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_46_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_46_io_wrEn = io_wrEn & io_wrTemplate == 7'h2e; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_46_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_46_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_47_clock = clock;
  assign templates_47_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_47_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_47_io_wrEn = io_wrEn & io_wrTemplate == 7'h2f; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_47_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_47_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_48_clock = clock;
  assign templates_48_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_48_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_48_io_wrEn = io_wrEn & io_wrTemplate == 7'h30; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_48_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_48_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_49_clock = clock;
  assign templates_49_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_49_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_49_io_wrEn = io_wrEn & io_wrTemplate == 7'h31; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_49_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_49_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_50_clock = clock;
  assign templates_50_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_50_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_50_io_wrEn = io_wrEn & io_wrTemplate == 7'h32; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_50_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_50_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_51_clock = clock;
  assign templates_51_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_51_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_51_io_wrEn = io_wrEn & io_wrTemplate == 7'h33; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_51_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_51_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_52_clock = clock;
  assign templates_52_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_52_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_52_io_wrEn = io_wrEn & io_wrTemplate == 7'h34; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_52_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_52_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_53_clock = clock;
  assign templates_53_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_53_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_53_io_wrEn = io_wrEn & io_wrTemplate == 7'h35; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_53_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_53_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_54_clock = clock;
  assign templates_54_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_54_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_54_io_wrEn = io_wrEn & io_wrTemplate == 7'h36; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_54_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_54_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_55_clock = clock;
  assign templates_55_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_55_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_55_io_wrEn = io_wrEn & io_wrTemplate == 7'h37; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_55_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_55_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_56_clock = clock;
  assign templates_56_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_56_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_56_io_wrEn = io_wrEn & io_wrTemplate == 7'h38; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_56_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_56_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_57_clock = clock;
  assign templates_57_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_57_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_57_io_wrEn = io_wrEn & io_wrTemplate == 7'h39; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_57_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_57_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_58_clock = clock;
  assign templates_58_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_58_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_58_io_wrEn = io_wrEn & io_wrTemplate == 7'h3a; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_58_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_58_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_59_clock = clock;
  assign templates_59_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_59_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_59_io_wrEn = io_wrEn & io_wrTemplate == 7'h3b; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_59_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_59_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_60_clock = clock;
  assign templates_60_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_60_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_60_io_wrEn = io_wrEn & io_wrTemplate == 7'h3c; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_60_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_60_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_61_clock = clock;
  assign templates_61_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_61_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_61_io_wrEn = io_wrEn & io_wrTemplate == 7'h3d; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_61_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_61_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_62_clock = clock;
  assign templates_62_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_62_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_62_io_wrEn = io_wrEn & io_wrTemplate == 7'h3e; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_62_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_62_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_63_clock = clock;
  assign templates_63_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_63_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_63_io_wrEn = io_wrEn & io_wrTemplate == 7'h3f; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_63_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_63_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_64_clock = clock;
  assign templates_64_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_64_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_64_io_wrEn = io_wrEn & io_wrTemplate == 7'h40; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_64_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_64_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_65_clock = clock;
  assign templates_65_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_65_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_65_io_wrEn = io_wrEn & io_wrTemplate == 7'h41; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_65_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_65_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_66_clock = clock;
  assign templates_66_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_66_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_66_io_wrEn = io_wrEn & io_wrTemplate == 7'h42; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_66_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_66_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_67_clock = clock;
  assign templates_67_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_67_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_67_io_wrEn = io_wrEn & io_wrTemplate == 7'h43; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_67_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_67_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_68_clock = clock;
  assign templates_68_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_68_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_68_io_wrEn = io_wrEn & io_wrTemplate == 7'h44; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_68_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_68_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_69_clock = clock;
  assign templates_69_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_69_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_69_io_wrEn = io_wrEn & io_wrTemplate == 7'h45; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_69_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_69_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_70_clock = clock;
  assign templates_70_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_70_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_70_io_wrEn = io_wrEn & io_wrTemplate == 7'h46; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_70_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_70_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_71_clock = clock;
  assign templates_71_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_71_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_71_io_wrEn = io_wrEn & io_wrTemplate == 7'h47; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_71_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_71_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_72_clock = clock;
  assign templates_72_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_72_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_72_io_wrEn = io_wrEn & io_wrTemplate == 7'h48; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_72_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_72_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_73_clock = clock;
  assign templates_73_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_73_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_73_io_wrEn = io_wrEn & io_wrTemplate == 7'h49; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_73_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_73_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_74_clock = clock;
  assign templates_74_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_74_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_74_io_wrEn = io_wrEn & io_wrTemplate == 7'h4a; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_74_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_74_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_75_clock = clock;
  assign templates_75_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_75_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_75_io_wrEn = io_wrEn & io_wrTemplate == 7'h4b; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_75_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_75_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_76_clock = clock;
  assign templates_76_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_76_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_76_io_wrEn = io_wrEn & io_wrTemplate == 7'h4c; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_76_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_76_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_77_clock = clock;
  assign templates_77_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_77_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_77_io_wrEn = io_wrEn & io_wrTemplate == 7'h4d; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_77_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_77_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_78_clock = clock;
  assign templates_78_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_78_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_78_io_wrEn = io_wrEn & io_wrTemplate == 7'h4e; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_78_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_78_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_79_clock = clock;
  assign templates_79_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_79_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_79_io_wrEn = io_wrEn & io_wrTemplate == 7'h4f; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_79_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_79_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_80_clock = clock;
  assign templates_80_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_80_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_80_io_wrEn = io_wrEn & io_wrTemplate == 7'h50; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_80_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_80_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_81_clock = clock;
  assign templates_81_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_81_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_81_io_wrEn = io_wrEn & io_wrTemplate == 7'h51; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_81_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_81_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_82_clock = clock;
  assign templates_82_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_82_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_82_io_wrEn = io_wrEn & io_wrTemplate == 7'h52; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_82_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_82_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_83_clock = clock;
  assign templates_83_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_83_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_83_io_wrEn = io_wrEn & io_wrTemplate == 7'h53; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_83_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_83_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_84_clock = clock;
  assign templates_84_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_84_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_84_io_wrEn = io_wrEn & io_wrTemplate == 7'h54; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_84_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_84_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_85_clock = clock;
  assign templates_85_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_85_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_85_io_wrEn = io_wrEn & io_wrTemplate == 7'h55; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_85_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_85_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_86_clock = clock;
  assign templates_86_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_86_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_86_io_wrEn = io_wrEn & io_wrTemplate == 7'h56; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_86_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_86_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_87_clock = clock;
  assign templates_87_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_87_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_87_io_wrEn = io_wrEn & io_wrTemplate == 7'h57; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_87_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_87_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_88_clock = clock;
  assign templates_88_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_88_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_88_io_wrEn = io_wrEn & io_wrTemplate == 7'h58; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_88_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_88_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_89_clock = clock;
  assign templates_89_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_89_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_89_io_wrEn = io_wrEn & io_wrTemplate == 7'h59; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_89_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_89_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_90_clock = clock;
  assign templates_90_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_90_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_90_io_wrEn = io_wrEn & io_wrTemplate == 7'h5a; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_90_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_90_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_91_clock = clock;
  assign templates_91_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_91_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_91_io_wrEn = io_wrEn & io_wrTemplate == 7'h5b; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_91_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_91_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_92_clock = clock;
  assign templates_92_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_92_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_92_io_wrEn = io_wrEn & io_wrTemplate == 7'h5c; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_92_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_92_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_93_clock = clock;
  assign templates_93_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_93_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_93_io_wrEn = io_wrEn & io_wrTemplate == 7'h5d; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_93_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_93_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_94_clock = clock;
  assign templates_94_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_94_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_94_io_wrEn = io_wrEn & io_wrTemplate == 7'h5e; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_94_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_94_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_95_clock = clock;
  assign templates_95_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_95_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_95_io_wrEn = io_wrEn & io_wrTemplate == 7'h5f; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_95_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_95_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_96_clock = clock;
  assign templates_96_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_96_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_96_io_wrEn = io_wrEn & io_wrTemplate == 7'h60; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_96_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_96_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_97_clock = clock;
  assign templates_97_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_97_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_97_io_wrEn = io_wrEn & io_wrTemplate == 7'h61; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_97_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_97_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_98_clock = clock;
  assign templates_98_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_98_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_98_io_wrEn = io_wrEn & io_wrTemplate == 7'h62; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_98_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_98_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
  assign templates_99_clock = clock;
  assign templates_99_io_lineAddr = io_lineAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 178:34]
  assign templates_99_io_lineEn = io_lineEn; // @[\\src\\main\\scala\\bram\\bramMem.scala 179:34]
  assign templates_99_io_wrEn = io_wrEn & io_wrTemplate == 7'h63; // @[\\src\\main\\scala\\bram\\bramMem.scala 183:43]
  assign templates_99_io_wrAddr = io_wrAddr; // @[\\src\\main\\scala\\bram\\bramMem.scala 184:32]
  assign templates_99_io_wrData = io_wrData; // @[\\src\\main\\scala\\bram\\bramMem.scala 185:32]
endmodule
